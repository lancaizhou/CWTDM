----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2018/04/20 16:14:54
-- Design Name: 
-- Module Name: synchronize - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity buhuo is
    Port ( clk_72M : in STD_LOGIC;
           data_in_i : in STD_LOGIC_VECTOR (15 downto 0);
		   data_in_q : in STD_LOGIC_VECTOR (15 downto 0);
			rst : in std_logic;
           sys_out : out STD_LOGIC_VECTOR (35 downto 0));
end buhuo;

architecture Behavioral of buhuo is
type tempp is array(511 downto 0) of std_logic_vector(17 downto 0);
signal xiangguan_i,xiangguan_q:tempp;
type Reg is array(511 downto 0) of std_logic_vector(15 downto 0);
signal regdin_i,regdin_q : Reg;
type PN_code is array(511 downto 0) of std_logic_vector(1 downto 0);
signal PN : PN_code:=("01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"00");
--先将I、Q两路信号相关

--相关峰
signal counter : std_logic_vector(14 downto 0);
--捕获使能信号
signal PN_en : std_logic;
signal dout_i : std_logic_vector(15 downto 0);
signal dout_q : std_logic_vector(15 downto 0);
begin
process(clk_72M,rst)
variable result_temp_i : std_logic_vector(17 downto 0);
variable result_temp_q : std_logic_vector(17 downto 0);
begin
	if rst='1' then
		regdin_i<=(others=>"0000000000000000");
		-- regdin_q<=(others=>"0000000000000000");
		regdin_q<=(others=>(others=>'0'));
		result_temp_i:=(others=>'0');
		result_temp_q:=(others=>'0');
		-- PN_en<='0';
		counter<=(others=>'0');
	elsif rising_edge(clk_72M) then
		for i in 0 to 511 loop
			if i=511 then
				regdin_i(i)<=data_in_i;
				regdin_q(i)<=data_in_q;
			else
				regdin_i(510-i)<=regdin_i(511-i);
				regdin_q(510-i)<=regdin_q(511-i);
			end if;
		end loop;
		
		-- for i in 0 to 511 loop
			-- regdin_i(i)<=xiangguan_i*PN(509-k);
		-- end loop;
		counter<=counter+1;
		result_temp_i:=(others=>'0');
		result_temp_q:=(others=>'0');
			for k in 0 to 510 loop
				result_temp_i:=result_temp_i+PN(510-k)*regdin_i(k);
				result_temp_q:=result_temp_q+PN(510-k)*regdin_q(k);
			end loop;	
			sys_out<=result_temp_i*result_temp_i+result_temp_q*result_temp_q;
			dout_i<=regdin_i(0);
			dout_q<=regdin_q(0);
	end if;
end process;
end Behavioral;








